module hello_world();

initial begin
	$display( "\n\tHello World!\n" );
end

endmodule
